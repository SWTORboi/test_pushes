module tonegen (
    input clk,
    input reset,
    input logic [7:0] volume,
    input logic [3:0] note,
    input logic [2:0] octave,
    input left_chan_ready,
    input right_chan_ready,
    output logic [15:0] sample_data,
    output logic sample_valid
);

		/* your code goes here */

endmodule